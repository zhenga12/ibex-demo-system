/* ------------------------------- 
 * RISC-V Vector LSU
 * ---------------------------------------------------------------------
 * Supporting:
 * VSEW: 8b, 16b, 32b
 * VLMUL: 1, 2, 4
 * Vector CSR:
 * 0x009    vxsat   fixed-point saturate flag
 * 0x00A    vxrm    fixed-point rounding mode (fixed to)
 * 0xC20    vl      vector length
 * 0xC21    vtype   vector data type register
 * 0xC22    vlenb   vector register length in bytes
 */
























